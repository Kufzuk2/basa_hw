
`define DISPLAY_0 7'b0111111
`define DISPLAY_OVERFLOW 7'b1100011

module numbers
(
    input   clk,
    input  KEY0, //reset
    input  KEY1, // translate
    input [7: 0] switches,

    output wire [7: 0] LEDR,
    output  reg [6: 0] HEX4, //right digit in hex
    output  reg [6: 0] HEX5, //left  digit in hex
    output  reg [6: 0] HEX6, //right digit in dec
    output  reg [6: 0] HEX7, //left  digit in dec

    output wire LEDG8
);

    assign LEDR = switches;

    // local hex ouputs
    wire [6: 0] hex4_loc;
    wire [6: 0] hex5_loc;
    wire [6: 0] hex6_loc;
    wire [6: 0] hex7_loc;
    

    wire [1: 0]    dec_offset;
    wire           dec_overflow; // might be replaced by ledg8
    assign LEDG8 = dec_overflow;


    // rst regs
    reg rst_push_1;
    reg rst_push_2;
    reg rst_pushed;

   
    // translate regs
    reg trans_push_1;
    reg trans_push_2;
    reg trans_pushed;


    // connection with decoder
    wire [3: 0]   hex_left;
    wire [3: 0]  hex_right;
    wire [3: 0]  dec_right;
    wire [3: 0]   dec_left;
    wire [7: 0] dec_in_hex;

    assign hex_left  =   switches[7: 4];
    assign hex_right =   switches[3: 0];
    assign dec_left  = dec_in_hex[7: 4];
    assign dec_right = dec_in_hex[3: 0];

    assign dec_overflow = (switches > 8'h63);

    decoder dec_hex_right
    (
        .HEX0(hex4_loc),
        .hex_num(hex_right)
    );

    decoder dec_hex_left
    (
        .HEX0(hex5_loc),
        .hex_num(hex_left)
    );

    decoder dec_dec_right
    (
        .HEX0(hex6_loc),
        .hex_num(dec_right)
    );

    decoder dec_dec_left
    (
        .HEX0(hex5_loc),
        .hex_num(dec_left)
    );


    // syncr reset logic
    always @(posedge clk) begin
        rst_push_1 <=       KEY0;
        rst_push_2 <= rst_push_1;
    end

    always @(posedge clk)
        rst_pushed <= ~rst_push_1 & rst_push_2;

        
    // syncr translation button logic
    always @(posedge clk) begin
        trans_push_1 <=         KEY0;
        trans_push_2 <= trans_push_1;
    end

    always @(posedge clk)
        trans_pushed <= ~trans_push_1 & trans_push_2;


    //hex display logic
    always @(posedge clk)
        if (rst_pushed) begin
            HEX4 <= `DISPLAY_0;  
            HEX5 <= `DISPLAY_0;  
        end else begin
            HEX4 <= trans_pushed ? hex4_loc : HEX4;  
            HEX5 <= trans_pushed ? hex5_loc : HEX5;  
        end


    //dec count logic
    genvar i;
    generate
        for (i = 0; i < 8; i = i + 1) begin
            if (i == 0) begin
                assign dec_in_hex = 0;
                assign dec_offset = 0;
            end else begin
                assign dec_in_hex = dec_in_hex + switches[i - 1] - (dec_in_hex > 8'h9) & 8'ha;
                assign dec_offset = dec_offset + (dec_in_hex > 9);
            end
        end
    endgenerate

    //dec display logic
    always @(posedge clk)
        if (rst_pushed) begin
            HEX6 <= `DISPLAY_0;  
            HEX7 <= `DISPLAY_0;  
        end else begin
            HEX6 <= ~trans_pushed ? HEX6 :
                     dec_overflow ? `DISPLAY_OVERFLOW : hex6_loc;  

            HEX7 <= ~trans_pushed ? HEX7 :
                     dec_overflow ? `DISPLAY_OVERFLOW : hex7_loc;  
        end

endmodule




