module decoder
(
    input  wire            clk,
    input  wire [3: 0] counter,
    output wire [6: 0]    HEX0
);



